module register_alias_table();

endmodule 