module reservation_station();

endmodule
