module instruction_buffer (equal, a, b); 


endmodule 