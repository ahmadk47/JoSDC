module mux2x1 #(parameter size = 32) (in1, in2, s, out);

	// inputs	
	input s;
	input [size - 1:0] in1, in2; // edited size
	
	// outputs
	output [size - 1:0] out;  // edited size

	// Unit logic
	assign out = (~s) ? in1 : in2;
	
endmodule