module common_data_bus();

endmodule 